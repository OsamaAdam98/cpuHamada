/* Team TECH GEEKS */
/*
*This file is to reduce the amount of magic numbers thrown in the code
*/
`define loadA 8'h00
`define loadB 8'h11
`define add 8'h2?
`define sub 8'h3?
`define multiply 8'h4?
`define divide 8'h5?
`define shiftLeft 8'h6?
`define shiftRight 8'h7?

//mode 1 constants

`define oneLoadA 8'h00
`define oneLoadB 8'h11
`define oneAdd 8'h22
`define oneSub 8'h33
`define oneMultiply 8'h44
`define oneDivide 8'h55
`define oneShiftLeft 8'h66
`define oneShiftRight 8'h77
