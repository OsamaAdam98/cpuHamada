/* Team TECH GEEKS */
/*
*This file is to reduce the amount of magic numbers thrown in the code
*/
`define loadA 8'h00
`define loadB 8'h11
`define add 8'h2?
`define sub 8'h3?
`define multiply 8'h4?
`define divide 8'h5?
`define shiftLeft 8'h6?
`define shiftRight 8'h7?